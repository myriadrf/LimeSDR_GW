// max10_onchipflash.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module max10_onchipflash (
		input  wire        clock,                   //    clk.clk
		input  wire        avmm_csr_addr,           //    csr.address
		input  wire        avmm_csr_read,           //       .read
		input  wire [31:0] avmm_csr_writedata,      //       .writedata
		input  wire        avmm_csr_write,          //       .write
		output wire [31:0] avmm_csr_readdata,       //       .readdata
		input  wire [17:0] avmm_data_addr,          //   data.address
		input  wire        avmm_data_read,          //       .read
		input  wire [31:0] avmm_data_writedata,     //       .writedata
		input  wire        avmm_data_write,         //       .write
		output wire [31:0] avmm_data_readdata,      //       .readdata
		output wire        avmm_data_waitrequest,   //       .waitrequest
		output wire        avmm_data_readdatavalid, //       .readdatavalid
		input  wire [3:0]  avmm_data_burstcount,    //       .burstcount
		input  wire        reset_n                  // nreset.reset_n
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       (""),
		.INIT_FILENAME_SIM                   (""),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M16SAU169I7G"),
		.DEVICE_ID                           ("16"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (4095),
		.SECTOR2_START_ADDR                  (4096),
		.SECTOR2_END_ADDR                    (8191),
		.SECTOR3_START_ADDR                  (8192),
		.SECTOR3_END_ADDR                    (47103),
		.SECTOR4_START_ADDR                  (47104),
		.SECTOR4_END_ADDR                    (75775),
		.SECTOR5_START_ADDR                  (75776),
		.SECTOR5_END_ADDR                    (143359),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (143359),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (8191),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (4),
		.SECTOR5_MAP                         (5),
		.ADDR_RANGE1_END_ADDR                (143359),
		.ADDR_RANGE2_END_ADDR                (143359),
		.ADDR_RANGE1_OFFSET                  (1024),
		.ADDR_RANGE2_OFFSET                  (0),
		.ADDR_RANGE3_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (18),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (4),
		.SECTOR_READ_PROTECTION_MODE         (0),
		.FLASH_SEQ_READ_DATA_COUNT           (4),
		.FLASH_ADDR_ALIGNMENT_BITS           (2),
		.FLASH_READ_CYCLE_MAX_INDEX          (4),
		.FLASH_RESET_CYCLE_MAX_INDEX         (20),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (96),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (28000000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (24400),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("True"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("True")
	) onchip_flash_0 (
		.clock                   (clock),                   //    clk.clk
		.reset_n                 (reset_n),                 // nreset.reset_n
		.avmm_data_addr          (avmm_data_addr),          //   data.address
		.avmm_data_read          (avmm_data_read),          //       .read
		.avmm_data_writedata     (avmm_data_writedata),     //       .writedata
		.avmm_data_write         (avmm_data_write),         //       .write
		.avmm_data_readdata      (avmm_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (avmm_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (avmm_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (avmm_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (avmm_csr_addr),           //    csr.address
		.avmm_csr_read           (avmm_csr_read),           //       .read
		.avmm_csr_writedata      (avmm_csr_writedata),      //       .writedata
		.avmm_csr_write          (avmm_csr_write),          //       .write
		.avmm_csr_readdata       (avmm_csr_readdata)        //       .readdata
	);

endmodule
